`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    03:03:08 11/10/2010 
// Design Name: 
// Module Name:    diff_select 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module diff_select( diff_p1p2, diff_p2p3, diff_p3p1, minp, diff_p1min, 
		    diff_p2minp, diff_p3minp);


endmodule
